// procesador.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module procesador (
		input  wire        clk_clk,                    //                  clk.clk
		output wire        enable_export,              //               enable.export
		input  wire        fifo_fft_imag_in_valid,     //     fifo_fft_imag_in.valid
		input  wire [31:0] fifo_fft_imag_in_data,      //                     .data
		input  wire        fifo_fft_real_in_valid,     //     fifo_fft_real_in.valid
		input  wire [31:0] fifo_fft_real_in_data,      //                     .data
		input  wire        fifo_resultados_cuad_valid, // fifo_resultados_cuad.valid
		input  wire [31:0] fifo_resultados_cuad_data,  //                     .data
		input  wire        fifo_resultados_fase_valid, // fifo_resultados_fase.valid
		input  wire [31:0] fifo_resultados_fase_data,  //                     .data
		output wire        pll_clock_clk,              //            pll_clock.clk
		input  wire        reset_reset_n,              //                reset.reset_n
		input  wire        reset_fifos_reset,          //          reset_fifos.reset
		output wire        reset_op_export             //             reset_op.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [18:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [18:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_resultados_fase_out_readdata;         // fifo_resultados_fase:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_resultados_fase_out_readdata
	wire   [0:0] mm_interconnect_0_fifo_resultados_fase_out_address;          // mm_interconnect_0:fifo_resultados_fase_out_address -> fifo_resultados_fase:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo_resultados_fase_out_read;             // mm_interconnect_0:fifo_resultados_fase_out_read -> fifo_resultados_fase:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_resultados_cuad_out_readdata;         // fifo_resultados_cuad:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_resultados_cuad_out_readdata
	wire   [0:0] mm_interconnect_0_fifo_resultados_cuad_out_address;          // mm_interconnect_0:fifo_resultados_cuad_out_address -> fifo_resultados_cuad:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo_resultados_cuad_out_read;             // mm_interconnect_0:fifo_resultados_cuad_out_read -> fifo_resultados_cuad:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_fft_real_out_readdata;                // fifo_fft_real:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_fft_real_out_readdata
	wire   [0:0] mm_interconnect_0_fifo_fft_real_out_address;                 // mm_interconnect_0:fifo_fft_real_out_address -> fifo_fft_real:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo_fft_real_out_read;                    // mm_interconnect_0:fifo_fft_real_out_read -> fifo_fft_real:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_fft_imag_out_readdata;                // fifo_fft_imag:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_fft_imag_out_readdata
	wire   [0:0] mm_interconnect_0_fifo_fft_imag_out_address;                 // mm_interconnect_0:fifo_fft_imag_out_address -> fifo_fft_imag:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo_fft_imag_out_read;                    // mm_interconnect_0:fifo_fft_imag_out_read -> fifo_fft_imag:avalonmm_read_slave_read
	wire         mm_interconnect_0_program_memory_s1_chipselect;              // mm_interconnect_0:program_memory_s1_chipselect -> program_memory:chipselect
	wire  [31:0] mm_interconnect_0_program_memory_s1_readdata;                // program_memory:readdata -> mm_interconnect_0:program_memory_s1_readdata
	wire  [14:0] mm_interconnect_0_program_memory_s1_address;                 // mm_interconnect_0:program_memory_s1_address -> program_memory:address
	wire   [3:0] mm_interconnect_0_program_memory_s1_byteenable;              // mm_interconnect_0:program_memory_s1_byteenable -> program_memory:byteenable
	wire         mm_interconnect_0_program_memory_s1_write;                   // mm_interconnect_0:program_memory_s1_write -> program_memory:write
	wire  [31:0] mm_interconnect_0_program_memory_s1_writedata;               // mm_interconnect_0:program_memory_s1_writedata -> program_memory:writedata
	wire         mm_interconnect_0_program_memory_s1_clken;                   // mm_interconnect_0:program_memory_s1_clken -> program_memory:clken
	wire         mm_interconnect_0_reset_s1_chipselect;                       // mm_interconnect_0:reset_s1_chipselect -> reset:chipselect
	wire  [31:0] mm_interconnect_0_reset_s1_readdata;                         // reset:readdata -> mm_interconnect_0:reset_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_s1_address;                          // mm_interconnect_0:reset_s1_address -> reset:address
	wire         mm_interconnect_0_reset_s1_write;                            // mm_interconnect_0:reset_s1_write -> reset:write_n
	wire  [31:0] mm_interconnect_0_reset_s1_writedata;                        // mm_interconnect_0:reset_s1_writedata -> reset:writedata
	wire         mm_interconnect_0_enable_s1_chipselect;                      // mm_interconnect_0:enable_s1_chipselect -> enable:chipselect
	wire  [31:0] mm_interconnect_0_enable_s1_readdata;                        // enable:readdata -> mm_interconnect_0:enable_s1_readdata
	wire   [1:0] mm_interconnect_0_enable_s1_address;                         // mm_interconnect_0:enable_s1_address -> enable:address
	wire         mm_interconnect_0_enable_s1_write;                           // mm_interconnect_0:enable_s1_write -> enable:write_n
	wire  [31:0] mm_interconnect_0_enable_s1_writedata;                       // mm_interconnect_0:enable_s1_writedata -> enable:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [enable:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, program_memory:reset, reset:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, program_memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [fifo_fft_imag:reset_n, fifo_fft_real:reset_n, fifo_resultados_cuad:reset_n, fifo_resultados_fase:reset_n, mm_interconnect_0:fifo_resultados_fase_reset_in_reset_bridge_in_reset_reset]

	procesador_enable enable (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_enable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_enable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_enable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_enable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_enable_s1_readdata),   //                    .readdata
		.out_port   (enable_export)                           // external_connection.export
	);

	procesador_fifo_fft_imag fifo_fft_imag (
		.wrclock                      (pll_clock_clk),                                //   clk_in.clk
		.reset_n                      (~rst_controller_001_reset_out_reset),          // reset_in.reset_n
		.avalonst_sink_valid          (fifo_fft_imag_in_valid),                       //       in.valid
		.avalonst_sink_data           (fifo_fft_imag_in_data),                        //         .data
		.avalonmm_read_slave_readdata (mm_interconnect_0_fifo_fft_imag_out_readdata), //      out.readdata
		.avalonmm_read_slave_read     (mm_interconnect_0_fifo_fft_imag_out_read),     //         .read
		.avalonmm_read_slave_address  (mm_interconnect_0_fifo_fft_imag_out_address)   //         .address
	);

	procesador_fifo_fft_imag fifo_fft_real (
		.wrclock                      (pll_clock_clk),                                //   clk_in.clk
		.reset_n                      (~rst_controller_001_reset_out_reset),          // reset_in.reset_n
		.avalonst_sink_valid          (fifo_fft_real_in_valid),                       //       in.valid
		.avalonst_sink_data           (fifo_fft_real_in_data),                        //         .data
		.avalonmm_read_slave_readdata (mm_interconnect_0_fifo_fft_real_out_readdata), //      out.readdata
		.avalonmm_read_slave_read     (mm_interconnect_0_fifo_fft_real_out_read),     //         .read
		.avalonmm_read_slave_address  (mm_interconnect_0_fifo_fft_real_out_address)   //         .address
	);

	procesador_fifo_resultados_cuad fifo_resultados_cuad (
		.wrclock                      (pll_clock_clk),                                       //   clk_in.clk
		.reset_n                      (~rst_controller_001_reset_out_reset),                 // reset_in.reset_n
		.avalonst_sink_valid          (fifo_resultados_cuad_valid),                          //       in.valid
		.avalonst_sink_data           (fifo_resultados_cuad_data),                           //         .data
		.avalonmm_read_slave_readdata (mm_interconnect_0_fifo_resultados_cuad_out_readdata), //      out.readdata
		.avalonmm_read_slave_read     (mm_interconnect_0_fifo_resultados_cuad_out_read),     //         .read
		.avalonmm_read_slave_address  (mm_interconnect_0_fifo_resultados_cuad_out_address)   //         .address
	);

	procesador_fifo_resultados_cuad fifo_resultados_fase (
		.wrclock                      (pll_clock_clk),                                       //   clk_in.clk
		.reset_n                      (~rst_controller_001_reset_out_reset),                 // reset_in.reset_n
		.avalonst_sink_valid          (fifo_resultados_fase_valid),                          //       in.valid
		.avalonst_sink_data           (fifo_resultados_fase_data),                           //         .data
		.avalonmm_read_slave_readdata (mm_interconnect_0_fifo_resultados_fase_out_readdata), //      out.readdata
		.avalonmm_read_slave_read     (mm_interconnect_0_fifo_resultados_fase_out_read),     //         .read
		.avalonmm_read_slave_address  (mm_interconnect_0_fifo_resultados_fase_out_address)   //         .address
	);

	procesador_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	procesador_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	procesador_pll_0 pll_0 (
		.refclk   (clk_clk),        //  refclk.clk
		.rst      (~reset_reset_n), //   reset.reset
		.outclk_0 (pll_clock_clk),  // outclk0.clk
		.locked   ()                // (terminated)
	);

	procesador_program_memory program_memory (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_program_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_program_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_program_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_program_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_program_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_program_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_program_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	procesador_enable reset (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_s1_readdata),   //                    .readdata
		.out_port   (reset_op_export)                        // external_connection.export
	);

	procesador_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                             (clk_clk),                                                     //                                           clk_0_clk.clk
		.pll_0_outclk0_clk                                         (pll_clock_clk),                                               //                                       pll_0_outclk0.clk
		.fifo_resultados_fase_reset_in_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // fifo_resultados_fase_reset_in_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                              //            nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                          (nios2_gen2_0_data_master_address),                            //                            nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                      (nios2_gen2_0_data_master_waitrequest),                        //                                                    .waitrequest
		.nios2_gen2_0_data_master_byteenable                       (nios2_gen2_0_data_master_byteenable),                         //                                                    .byteenable
		.nios2_gen2_0_data_master_read                             (nios2_gen2_0_data_master_read),                               //                                                    .read
		.nios2_gen2_0_data_master_readdata                         (nios2_gen2_0_data_master_readdata),                           //                                                    .readdata
		.nios2_gen2_0_data_master_write                            (nios2_gen2_0_data_master_write),                              //                                                    .write
		.nios2_gen2_0_data_master_writedata                        (nios2_gen2_0_data_master_writedata),                          //                                                    .writedata
		.nios2_gen2_0_data_master_debugaccess                      (nios2_gen2_0_data_master_debugaccess),                        //                                                    .debugaccess
		.nios2_gen2_0_instruction_master_address                   (nios2_gen2_0_instruction_master_address),                     //                     nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest               (nios2_gen2_0_instruction_master_waitrequest),                 //                                                    .waitrequest
		.nios2_gen2_0_instruction_master_read                      (nios2_gen2_0_instruction_master_read),                        //                                                    .read
		.nios2_gen2_0_instruction_master_readdata                  (nios2_gen2_0_instruction_master_readdata),                    //                                                    .readdata
		.enable_s1_address                                         (mm_interconnect_0_enable_s1_address),                         //                                           enable_s1.address
		.enable_s1_write                                           (mm_interconnect_0_enable_s1_write),                           //                                                    .write
		.enable_s1_readdata                                        (mm_interconnect_0_enable_s1_readdata),                        //                                                    .readdata
		.enable_s1_writedata                                       (mm_interconnect_0_enable_s1_writedata),                       //                                                    .writedata
		.enable_s1_chipselect                                      (mm_interconnect_0_enable_s1_chipselect),                      //                                                    .chipselect
		.fifo_fft_imag_out_address                                 (mm_interconnect_0_fifo_fft_imag_out_address),                 //                                   fifo_fft_imag_out.address
		.fifo_fft_imag_out_read                                    (mm_interconnect_0_fifo_fft_imag_out_read),                    //                                                    .read
		.fifo_fft_imag_out_readdata                                (mm_interconnect_0_fifo_fft_imag_out_readdata),                //                                                    .readdata
		.fifo_fft_real_out_address                                 (mm_interconnect_0_fifo_fft_real_out_address),                 //                                   fifo_fft_real_out.address
		.fifo_fft_real_out_read                                    (mm_interconnect_0_fifo_fft_real_out_read),                    //                                                    .read
		.fifo_fft_real_out_readdata                                (mm_interconnect_0_fifo_fft_real_out_readdata),                //                                                    .readdata
		.fifo_resultados_cuad_out_address                          (mm_interconnect_0_fifo_resultados_cuad_out_address),          //                            fifo_resultados_cuad_out.address
		.fifo_resultados_cuad_out_read                             (mm_interconnect_0_fifo_resultados_cuad_out_read),             //                                                    .read
		.fifo_resultados_cuad_out_readdata                         (mm_interconnect_0_fifo_resultados_cuad_out_readdata),         //                                                    .readdata
		.fifo_resultados_fase_out_address                          (mm_interconnect_0_fifo_resultados_fase_out_address),          //                            fifo_resultados_fase_out.address
		.fifo_resultados_fase_out_read                             (mm_interconnect_0_fifo_resultados_fase_out_read),             //                                                    .read
		.fifo_resultados_fase_out_readdata                         (mm_interconnect_0_fifo_resultados_fase_out_readdata),         //                                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_address                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                    .write
		.jtag_uart_0_avalon_jtag_slave_read                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                    .chipselect
		.nios2_gen2_0_debug_mem_slave_address                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //                        nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                                    .write
		.nios2_gen2_0_debug_mem_slave_read                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                                    .read
		.nios2_gen2_0_debug_mem_slave_readdata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                                    .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                                    .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                                    .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                                    .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                                    .debugaccess
		.program_memory_s1_address                                 (mm_interconnect_0_program_memory_s1_address),                 //                                   program_memory_s1.address
		.program_memory_s1_write                                   (mm_interconnect_0_program_memory_s1_write),                   //                                                    .write
		.program_memory_s1_readdata                                (mm_interconnect_0_program_memory_s1_readdata),                //                                                    .readdata
		.program_memory_s1_writedata                               (mm_interconnect_0_program_memory_s1_writedata),               //                                                    .writedata
		.program_memory_s1_byteenable                              (mm_interconnect_0_program_memory_s1_byteenable),              //                                                    .byteenable
		.program_memory_s1_chipselect                              (mm_interconnect_0_program_memory_s1_chipselect),              //                                                    .chipselect
		.program_memory_s1_clken                                   (mm_interconnect_0_program_memory_s1_clken),                   //                                                    .clken
		.reset_s1_address                                          (mm_interconnect_0_reset_s1_address),                          //                                            reset_s1.address
		.reset_s1_write                                            (mm_interconnect_0_reset_s1_write),                            //                                                    .write
		.reset_s1_readdata                                         (mm_interconnect_0_reset_s1_readdata),                         //                                                    .readdata
		.reset_s1_writedata                                        (mm_interconnect_0_reset_s1_writedata),                        //                                                    .writedata
		.reset_s1_chipselect                                       (mm_interconnect_0_reset_s1_chipselect)                        //                                                    .chipselect
	);

	procesador_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (reset_fifos_reset),                  // reset_in1.reset
		.clk            (pll_clock_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
